// ============================================================================
// Copyright (c) 2016 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//  
//  
//                     web: http://www.terasic.com/  
//                     email: support@terasic.com
//
// ============================================================================
//Date:  Wed May 11 09:51:57 2016
// ============================================================================

module DE10_LITE_GSensor(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// VGA //////////
	output		     [3:0]		VGA_B,
	output		     [3:0]		VGA_G,
	output		          		VGA_HS,
	output		     [3:0]		VGA_R,
	output		          		VGA_VS,

	//////////// Accelerometer //////////
	output		          		GSENSOR_CS_N,
	input 		     [2:1]		GSENSOR_INT,
	output		          		GSENSOR_SCLK,
	output		          		GSENSOR_SDI,
	input 		          		GSENSOR_SDO,

	//////////// Arduino //////////
	inout 		    [15:0]		ARDUINO_IO,
	inout 		          		ARDUINO_RESET_N,
	///////HEX//////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4
);

//=======================================================
//  REG/WIRE declarations
//=======================================================
wire	        dly_rst;
wire	        spi_clk, spi_clk_out;
wire	[15:0]  data_x;
wire	[15:0]  data_y;
//=======================================================
//  7-segment 지연 출력 wire / reg
//=======================================================
wire [6:0]hex0;
wire [6:0]hex1;
wire [6:0]hex2;
wire [6:0]hex3;
wire[6:0]hex4;

reg[6:0]h0;
reg[6:0]h1;
reg[6:0]h2;
reg[6:0]h3;
reg[6:0]h4;

reg [25:0] count;


//=======================================================
//  Structural coding
//=======================================================

//	Reset
reset_delay	u_reset_delay	(	
            .iRSTN(KEY[1]),
            .iCLK(MAX10_CLK1_50),
            .oRST(dly_rst));

//  PLL            
spi_pll     u_spi_pll	(
            .areset(dly_rst),
            .inclk0(MAX10_CLK1_50),
            .c0(spi_clk),      // 2MHz
            .c1(spi_clk_out)); // 2MHz phase shift 

//  Initial Setting and Data Read Back
spi_ee_config u_spi_ee_config (			
						.iRSTN(!dly_rst),															
						.iSPI_CLK(spi_clk),								
						.iSPI_CLK_OUT(spi_clk_out),								
						.iG_INT2(GSENSOR_INT[1]),            
						.oDATA_L(data_x[7:0]),
						.oDATA_H(data_x[15:8]),
						.oY_DATA_L(data_y[7:0]),
						.oY_DATA_H(data_y[15:8]),
						.oSPI_SDI(GSENSOR_SDI),
						.iSPI_SDO(GSENSOR_SDO),
						.oSPI_CSN(GSENSOR_CS_N),
						.oSPI_CLK(GSENSOR_SCLK),
						.HEX0(hex0),
						.HEX1(hex1),
						.HEX2(hex2),
						.HEX3(hex3),
						.HEX4(hex4));
			
//	LED
led_driver u_led_driver	(	
						.iRSTN(!dly_rst),
						.iCLK(MAX10_CLK1_50),
						.iDIG(data_x[9:0]),
						.iG_INT2(GSENSOR_INT[1]),            
						.oLED(LEDR));

// VGA: black background with white dot controlled by X/Y tilt
vga_tilt_dot u_vga_tilt_dot(
						.iCLK(MAX10_CLK1_50),
						.iRST(dly_rst),
						.iDRAW_EN(!KEY[0]),
						.iTILT_X(data_x),
						.iTILT_Y(data_y),
						.oVGA_R(VGA_R),
						.oVGA_G(VGA_G),
						.oVGA_B(VGA_B),
						.oVGA_HS(VGA_HS),
						.oVGA_VS(VGA_VS));

// 1초 지연을 위한 카운터
always@(posedge MAX10_CLK1_50 or posedge dly_rst)
begin
	if (dly_rst)
	begin
		count <= 1'b0;
	end
	else
	begin
		
		if (count==26'd50_000_000) // 1초 지연
		begin
			count <= 1'b0;
			h0 <= hex0;
			h1 <= hex1;
			h2 <= hex2;
			h3 <= hex3;
			h4 <= hex4;
		end
		else
		begin
			count <= count+1'b1;
			h0 <= h0;
			h1 <= h1;
			h2 <= h2;
			h3 <= h3;
			h4 <= h4;
		end
	end
end

assign HEX0 = h0;
assign HEX1 = h1;
assign HEX2 = h2;
assign HEX3 = h3;
assign HEX4 = h4;



endmodule
